module SidewalkLight(clk,rows,cols);
input clk;
output reg [15:0] rows;
output reg [3:0] cols;

reg [4:0] state;
reg [9:0] cnt;
reg walk;

always @(posedge clk) begin
	 cnt=cnt+1;
	 cols=cols+1;
	 
	 if(cnt==10'b1111111111) begin
	     cnt=10'b0000000000;
		  walk=~walk;
	 end
	 
end

always @(cnt[5]) begin
   state=state+1;
	if(walk) begin
	     if(state==5'b10001) state=5'b00000;
	 end
	 else begin
	     state=5'b10010;
	 end
end

always @(cols) begin
    if(state==5'b00000) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000010000100;
				4: rows=16'b0111000100000100;
				5: rows=16'b0111111100001000;
				6: rows=16'b0010111100010000;
				7: rows=16'b0000011111100000;
				8: rows=16'b0000010011000000;
				9: rows=16'b0000001000100000;
				10: rows=16'b0000000000010000;
				11: rows=16'b0000000000001000;
				12: rows=16'b0000000000000110;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b0001) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000010000110;
				4: rows=16'b0111000110000110;
				5: rows=16'b0111111100001010;
				6: rows=16'b0010111100011100;
				7: rows=16'b0000011111100000;
				8: rows=16'b0000010011000000;
				9: rows=16'b0000011000100000;
				10: rows=16'b0000001110010010;
				11: rows=16'b0000000100011010;
				12: rows=16'b0000000000001110;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b00010) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000000000010;
				4: rows=16'b0111000010000010;
				5: rows=16'b0111111100000010;
				6: rows=16'b0010111100011100;
				7: rows=16'b0000011111100000;
				8: rows=16'b0000010011000000;
				9: rows=16'b0000010000100000;
				10: rows=16'b0000001000010000;
				11: rows=16'b0000000100010010;
				12: rows=16'b0000000000001100;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b00011) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000000000000;
				4: rows=16'b0111000010000010;
				5: rows=16'b0111111100011010;
				6: rows=16'b0010111100100110;
				7: rows=16'b0000010111000000;
				8: rows=16'b0000010011000000;
				9: rows=16'b0000001000110100;
				10: rows=16'b0000000110010100;
				11: rows=16'b0000000000011000;
				12: rows=16'b0000000000000000;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b00100) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000000000000;
				4: rows=16'b0111000010000010;
				5: rows=16'b0111111100011111;
				6: rows=16'b0010111110100111;
				7: rows=16'b0000010111100000;
				8: rows=16'b0000011011110000;
				9: rows=16'b0000001110111100;
				10: rows=16'b0000000110011100;
				11: rows=16'b0000000000011110;
				12: rows=16'b0000000000000000;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b00101) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000000000000;
				4: rows=16'b0111000000000000;
				5: rows=16'b0111111000010101;
				6: rows=16'b0010111110100111;
				7: rows=16'b0000010111100000;
				8: rows=16'b0000001001110000;
				9: rows=16'b0000000110001000;
				10: rows=16'b0000000000001000;
				11: rows=16'b0000000000000110;
				12: rows=16'b0000000000000000;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b00110) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000000000000;
				4: rows=16'b0111000000011001;
				5: rows=16'b0111111010100101;
				6: rows=16'b0010111111100111;
				7: rows=16'b0000010111110000;
				8: rows=16'b0000001000001000;
				9: rows=16'b0000000000000110;
				10: rows=16'b0000000000000000;
				11: rows=16'b0000000000000000;
				12: rows=16'b0000000000000000;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b00111) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000000000000;
				4: rows=16'b0111000000000000;
				5: rows=16'b0111111000100000;
				6: rows=16'b0010111111000000;
				7: rows=16'b0000011111111010;
				8: rows=16'b0000000011101000;
				9: rows=16'b0000000000111110;
				10: rows=16'b0000000000000000;
				11: rows=16'b0000000000000000;
				12: rows=16'b0000000000000000;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b01000) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000000000000;
				4: rows=16'b0111000100000100;
				5: rows=16'b0111110100010100;
				6: rows=16'b0010111111101100;
				7: rows=16'b0000011111110000;
				8: rows=16'b0000011111111010;
				9: rows=16'b0000001100001001;
				10: rows=16'b0000000000000111;
				11: rows=16'b0000000000000001;
				12: rows=16'b0000000000000000;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b01001) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000000000000;
				4: rows=16'b0111000000000000;
				5: rows=16'b0111111000010101;
				6: rows=16'b0010111110100111;
				7: rows=16'b0000011111110000;
				8: rows=16'b0000011111111010;
				9: rows=16'b0000001100001001;
				10: rows=16'b0000000000000111;
				11: rows=16'b0000000000000001;
				12: rows=16'b0000000000000000;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b01010) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000000000001;
				4: rows=16'b0111000010000001;
				5: rows=16'b0111111100000001;
				6: rows=16'b0010111100011110;
				7: rows=16'b0000011111100000;
				8: rows=16'b0000010011000000;
				9: rows=16'b0000010000100000;
				10: rows=16'b0000001000010000;
				11: rows=16'b0000000100010010;
				12: rows=16'b0000000000001100;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b01011) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000000000000;
				4: rows=16'b0111000010000010;
				5: rows=16'b0111111100011010;
				6: rows=16'b0010111100100110;
				7: rows=16'b0000010111000000;
				8: rows=16'b0000010011000000;
				9: rows=16'b0000001000110100;
				10: rows=16'b0000000110010100;
				11: rows=16'b0000000000011000;
				12: rows=16'b0000000000000000;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b01100) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000000000000;
				4: rows=16'b0111111000011101;
				5: rows=16'b0111111110100111;
				6: rows=16'b0010111111100111;
				7: rows=16'b0000011111110000;
				8: rows=16'b0000001110001000;
				9: rows=16'b0000000000001110;
				10: rows=16'b0000000000000110;
				11: rows=16'b0000000000000000;
				12: rows=16'b0000000000000000;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b01101) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000000000000;
				4: rows=16'b0111000000011001;
				5: rows=16'b0111111010100101;
				6: rows=16'b0010111111100111;
				7: rows=16'b0000010111110000;
				8: rows=16'b0000001000001000;
				9: rows=16'b0000000000000110;
				10: rows=16'b0000000000000000;
				11: rows=16'b0000000000000000;
				12: rows=16'b0000000000000000;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b01110) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000000000000;
				4: rows=16'b0111000000000000;
				5: rows=16'b0111111000100000;
				6: rows=16'b0010111111000000;
				7: rows=16'b0000011111111010;
				8: rows=16'b0000000011101000;
				9: rows=16'b0000000000111110;
				10: rows=16'b0000000000000000;
				11: rows=16'b0000000000000000;
				12: rows=16'b0000000000000000;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b01111) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000000000000;
				4: rows=16'b0111000100000100;
				5: rows=16'b0111110100010100;
				6: rows=16'b0010111111101100;
				7: rows=16'b0000011111110000;
				8: rows=16'b0000011111111010;
				9: rows=16'b0000001100001001;
				10: rows=16'b0000000000000111;
				11: rows=16'b0000000000000001;
				12: rows=16'b0000000000000000;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b10000) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000010000100;
				4: rows=16'b0111000100000100;
				5: rows=16'b0111111100011100;
				6: rows=16'b0010111111111100;
				7: rows=16'b0000011111110000;
				8: rows=16'b0000011111111010;
				9: rows=16'b0000001100101001;
				10: rows=16'b0000000110010111;
				11: rows=16'b0000000000001001;
				12: rows=16'b0000000000000110;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b10001) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0010000010000100;
				4: rows=16'b0111000100000100;
				5: rows=16'b0111111100001000;
				6: rows=16'b0010111100010000;
				7: rows=16'b0000011111100000;
				8: rows=16'b0000011111100000;
				9: rows=16'b0000001000100000;
				10: rows=16'b0000000110010000;
				11: rows=16'b0000000000001000;
				12: rows=16'b0000000000000110;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
	 if(state==5'b10010) begin
	     case(cols)
		      0: rows=16'b0000000000000000;
				1: rows=16'b0000000000000000;
				2: rows=16'b0000000000000000;
				3: rows=16'b0000000000000000;
				4: rows=16'b0000001111110011;
				5: rows=16'b0000011111100011;
				6: rows=16'b0000111100011111;
				7: rows=16'b0111111111111111;
				8: rows=16'b0111111111110000;
				9: rows=16'b0111111111111111;
				10: rows=16'b0000111100011111;
				11: rows=16'b0000011111100011;
				12: rows=16'b0000001111110011;
				13: rows=16'b0000000000000000;
				14: rows=16'b0000000000000000;
				15: rows=16'b0000000000000000;
		  endcase
	 end
end

endmodule